// constraint constraint_identifier {variable dist{set of legal values and weights};}
