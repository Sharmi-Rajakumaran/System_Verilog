class enc;
  mailbox #(trans) gen2drv = new();
  
