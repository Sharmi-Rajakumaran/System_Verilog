// pattern 021346578







// pattern 0102030405
