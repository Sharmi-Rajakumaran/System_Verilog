class parent;
  rand bit [2:0]a;
  constraint a_size {a == 3;}
endclass: parent
